library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;

library work;
use work.TdmaMinTypes.all;

entity AVGASP_Wave_Test is
    generic (
        ports : positive := 8
    );
end entity;

architecture sim of AVGASP_Wave_Test is
    signal clock: STD_LOGIC:='1';
    signal send_port : tdma_min_ports(0 to ports-1);
    signal recv_port : tdma_min_ports(0 to ports-1);
    signal flag: STD_LOGIC:='0';

begin

    clock<= not clock after 10 ns;
    flag<= '1' after 50 ns;
	 
	 
    tdma_min: entity work.TdmaMin
        generic map (
            ports => ports
        )
        port map (
            clock => clock,
            sends => send_port,
            recvs => recv_port
        );

    avgCalc_ASP: entity work.AverageCalculator
        port map(
             clk    => clock,
				 reset  => '0',
		  
				 recv   => recv_port(2),  	  
		       send	  => send_port(2)
        );

--     test_Config: entity work.TestConfig
--        port map(
--			  clock => clock,
--			  send  => send_port(1),
--			  recv  => recv_port(1),
--			  flag => flag
--        );
		  
      test_ADC: entity work.TestAdc
	generic map(
		forward => 2
		)
        port map(
			  flag => flag,
			  clock => clock,
			  send  => send_port(0),
			  recv  => recv_port(0)
        );
	 
end architecture;